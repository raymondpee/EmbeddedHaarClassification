module database_embedded
#(
parameter ADDR_WIDTH = 10,
parameter DATA_WIDTH_8 = 8,   
parameter DATA_WIDTH_12 = 12, 
parameter DATA_WIDTH_16 = 16, 
parameter NUM_PARAM_PER_CLASSIFIER= 19,
parameter NUM_STAGE_THRESHOLD = 3,
parameter FILE_STAGE_FILE_1 = "memory1.mif",
parameter FILE_STAGE_FILE_2 = "memory2.mif",
parameter FILE_STAGE_FILE_3 = "memory3.mif",
parameter NUM_CLASSIFIERS_STAGE_1 = 10,
parameter NUM_CLASSIFIERS_STAGE_2 = 10,
parameter NUM_CLASSIFIERS_STAGE_3 = 10
)
(
clk,
reset,

)

input clk;
input reset;
output [DATA_WIDTH_16-1:0] o_memory[TOTAL_SIZE-1:0];


localparam SIZE_STAGE_1 = NUM_CLASSIFIERS_STAGE_1*NUM_PARAM_PER_CLASSIFIER + NUM_STAGE_THRESHOLD;
localparam SIZE_STAGE_2 = NUM_CLASSIFIERS_STAGE_2*NUM_PARAM_PER_CLASSIFIER + NUM_STAGE_THRESHOLD;
localparam SIZE_STAGE_3 = NUM_CLASSIFIERS_STAGE_3*NUM_PARAM_PER_CLASSIFIER + NUM_STAGE_THRESHOLD;
localparam TOTAL_SIZE = SIZE_STAGE_1 + SIZE_STAGE_2 + SIZE_STAGE_3;

reg[DATA_WIDTH_16-1:0] memory[TOTAL_SIZE-1:0];



assign o_memory = memory;


database_stage_memory
#(
.ADDR_WIDTH(ADDR_WIDTH),
.FILE_STAGE_MEM(FILE_STAGE_MEM),
.SIZE_STAGE(SIZE_STAGE)
)
database_stage_memory
(
.clk(clk),
.reset(reset),
.ren_database_index(renable),
.ren_database(renable),
.o_data(data)
);

endmodule